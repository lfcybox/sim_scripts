**.subckt test_sch
V1 IN GND pulse 0 3 '0.495/ 10e6 ' '0.01/10e6 ' '0.01/10e6 ' '0.49/10e6 ' '1/10e6 ' 
R1 OUT IN 100k m=1
R2 GND OUT 100k m=1
C1 OUT GND 10p m=1
**** begin user architecture code


.save all
.tran 1n 1u
.plot IN OUT


**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.end
